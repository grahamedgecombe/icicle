// Defines for Upduino
`define FLASH

