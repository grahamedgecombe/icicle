`ifndef RV32_MEM_OPS
`define RV32_MEM_OPS

localparam RV32_MEM_WIDTH_WORD = 2'b00;
localparam RV32_MEM_WIDTH_HALF = 2'b01;
localparam RV32_MEM_WIDTH_BYTE = 2'b10;

`endif
