// Defines for Icebreaker
`define SPI_FLASH
`define INTERNAL_OSC
