// Defines for BlackIce-II

