// Defines for iCE40-HX8K breakout board
//`define SPI_FLASH
