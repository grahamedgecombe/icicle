// Defines for Upduino
`define FLASH
`define INTERNAL_OSC
