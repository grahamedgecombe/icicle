module pll (
    input clock_in,
    output logic clock_out,
    output logic locked
);
    EHXPLLL #(
        .PLLRST_ENA("DISABLED"),
        .INTFB_WAKE("DISABLED"),
        .STDBY_ENABLE("DISABLED"),
        .DPHASE_SOURCE("DISABLED"),
        .CLKOS3_FPHASE(0),
        .CLKOS3_CPHASE(0),
        .CLKOS2_FPHASE(0),
        .CLKOS2_CPHASE(0),
        .CLKOS_FPHASE(0),
        .CLKOS_CPHASE(0),
        .CLKOP_FPHASE(0),
        .CLKOP_CPHASE(11),
        .PLL_LOCK_MODE(0),
        .CLKOS_TRIM_DELAY(0),
        .CLKOS_TRIM_POL("FALLING"),
        .CLKOP_TRIM_DELAY(0),
        .CLKOP_TRIM_POL("FALLING"),
        .OUTDIVIDER_MUXD("DIVD"),
        .CLKOS3_ENABLE("DISABLED"),
        .OUTDIVIDER_MUXC("DIVC"),
        .CLKOS2_ENABLE("DISABLED"),
        .OUTDIVIDER_MUXB("DIVB"),
        .CLKOS_ENABLE("DISABLED"),
        .OUTDIVIDER_MUXA("DIVA"),
        .CLKOP_ENABLE("ENABLED"),
        .CLKOS3_DIV(1),
        .CLKOS2_DIV(1),
        .CLKOS_DIV(1),
        .CLKOP_DIV(12),
        .CLKFB_DIV(4),
        .CLKI_DIV(1),
        .FEEDBK_PATH("CLKOP")
    ) pll (
        .CLKI(clock_in),
        .CLKFB(clock_out),
        .PHASESEL1(0),
        .PHASESEL0(0),
        .PHASEDIR(0),
        .PHASESTEP(0),
        .PHASELOADREG(0),
        .STDBY(0),
        .PLLWAKESYNC(0),
        .RST(0),
        .ENCLKOP(0),
        .ENCLKOS(0),
        .ENCLKOS2(0),
        .ENCLKOS3(0),
        .CLKOP(clock_out),
        .LOCK(locked)
    );
endmodule
